module HLSM (Clk, Rst, Start, Done);
	input Clk, Rst, Start;
	output reg Done;
	
	always @(posedge Clk) begin
			
	end
	
endmodule